`default_nettype none
module decoder_sim
  (input wire        wb_clk,
   input wire [31:2] wb_rdt,
   input wire        wb_en,
   output wire       ebreak,
   output wire       jal_or_jalr,
   output wire       mret,
   output wire       wfi,
   output wire       sh_right,
   output wire       bne_or_bge,
   output wire       cond_branch,
   output wire       e_op,
   output wire       branch_op,
   output wire       shift_op,
   output wire       slt_or_branch,
   output wire       rd_op,
   output wire       two_stage_op,
   output wire       dbus_en,
   output wire       mdu_op,
   output wire [2:0] ext_funct3,
   output wire       bufreg_rs1_en,
   output wire       bufreg_imm_en,
   output wire       bufreg_clr_lsb,
   output wire       bufreg_sh_signed,
   output wire       ctrl_utype,
   output wire       ctrl_pc_rel,
   output wire       alu_sub,
   output wire [1:0] alu_bool_op,
   output wire       alu_cmp_eq,
   output wire       alu_cmp_sig,
   output wire [2:0] alu_rd_sel,
   output wire       mem_signed,
   output wire       mem_word,
   output wire       mem_half,
   output wire       mem_cmd,
   output wire       csr_en,
   output wire [1:0] csr_addr,
   output wire       csr_mstatus_en,
   output wire       csr_mie_en,
   output wire       csr_mcause_en,
   output wire [1:0] csr_source,
   output wire       csr_d_sel,
   output wire       csr_imm_en,
   output wire       mtval_pc,
   output wire [3:0] immdec_ctrl,
   output wire [3:0] immdec_en,
   output wire       op_b_source,
   output wire       rd_mem_en,
   output wire       rd_csr_en,
   output wire       rd_alu_en
);

   // Instantiate the DUT
   serv_decode
     #(.PRE_REGISTER (1),
       .MDU (0))
   dut (
       .clk(wb_clk),
       .i_wb_rdt(wb_rdt),
       .i_wb_en(wb_en),
       // Outputs
       .o_sh_right(sh_right),
       .o_bne_or_bge(bne_or_bge),
       .o_cond_branch(cond_branch),
       .o_e_op(e_op),
       .o_ebreak(ebreak),
       .o_wfi(wfi),
       .o_branch_op(branch_op),
       .o_shift_op(shift_op),
       .o_slt_or_branch(slt_or_branch),
       .o_rd_op(rd_op),
       .o_two_stage_op(two_stage_op),
       .o_dbus_en(dbus_en),
       .o_mdu_op(mdu_op),
       .o_ext_funct3(ext_funct3),
       .o_bufreg_rs1_en(bufreg_rs1_en),
       .o_bufreg_imm_en(bufreg_imm_en),
       .o_bufreg_clr_lsb(bufreg_clr_lsb),
       .o_bufreg_sh_signed(bufreg_sh_signed),
       .o_ctrl_jal_or_jalr(jal_or_jalr),
       .o_ctrl_utype(ctrl_utype),
       .o_ctrl_pc_rel(ctrl_pc_rel),
       .o_ctrl_mret(mret),
       .o_alu_sub(alu_sub),
       .o_alu_bool_op(alu_bool_op),
       .o_alu_cmp_eq(alu_cmp_eq),
       .o_alu_cmp_sig(alu_cmp_sig),
       .o_alu_rd_sel(alu_rd_sel),
       .o_mem_signed(mem_signed),
       .o_mem_word(mem_word),
       .o_mem_half(mem_half),
       .o_mem_cmd(mem_cmd),
       .o_csr_en(csr_en),
       .o_csr_addr(csr_addr),
       .o_csr_mstatus_en(csr_mstatus_en),
       .o_csr_mie_en(csr_mie_en),
       .o_csr_mcause_en(csr_mcause_en),
       .o_csr_source(csr_source),
       .o_csr_d_sel(csr_d_sel),
       .o_csr_imm_en(csr_imm_en),
       .o_mtval_pc(mtval_pc),
       .o_immdec_ctrl(immdec_ctrl),
       .o_immdec_en(immdec_en),
       .o_op_b_source(op_b_source),
       .o_rd_mem_en(rd_mem_en),
       .o_rd_csr_en(rd_csr_en),
       .o_rd_alu_en(rd_alu_en)
   );

endmodule
